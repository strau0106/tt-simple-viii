package control;
    typedef enum {LEFT, RIGHT} op_dir_e /*verilator public*/;
    typedef enum {ADD, SUB, MUL, DIV, SHIFTL, ROTL, SHIFTR, ROTR, AND, OR, XOR, NOT} alu_op_e /*verilator public*/;
endpackage
