package control;
    typedef enum {LEFT, RIGHT} op_dir_e /*verilator public*/;
endpackage